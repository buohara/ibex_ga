// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * GA-Extended Ibex ID Stage
 * 
 * This module extends the original ibex_id_stage with GA coprocessor integration.
 * For now this is a placeholder that includes the original ID stage.
 */

// For now, just include the original ibex_id_stage  
// This will be extended later with actual GA integration
`include "../../../rtl/ibex_id_stage.sv"
